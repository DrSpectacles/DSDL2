module dot_adder(input [6:0] pattern,
		 
		 );
   
